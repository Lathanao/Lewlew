module classes

//import crypto.sha256
//import rand
//import os
//import time
//import sqlite

struct AdminFactory {
}
