// Copyright (c) 2019-2020 Alexander Medvednikov. All rights reserved.
// Use of this source code is governed by a GPL license that can be found in the LICENSE file.
module classes

struct Admin {
	AdminAbstract
	AdminFilter
	AdminEntity
}