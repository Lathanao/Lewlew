module dashboard
