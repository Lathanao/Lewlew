module classes

pub struct Tool {
}

pub fn (t Tool) display_error(error string, htmlentities bool) string {
	// global $_ERRORS;

	// if (is_null($context)) {
	// 		$context = Context::getContext();
	// }

	// @include_once(_PS_TRANSLATIONS_DIR_.$context->language->iso_code.'/errors.php');

	// if (defined('_PS_MODE_DEV_') && _PS_MODE_DEV_ && $string == 'Fatal error') {
	// 		return ('<pre>'.print_r(debug_backtrace(), true).'</pre>');
	// }

	// $key = md5(str_replace('\'', '\\\'', $string));
	// if (isset($_ERRORS)
	// 		&& is_array($_ERRORS)
	// 		&& array_key_exists($key, $_ERRORS)
	// 		&& $_ERRORS[$key] !== '') {
	// 		$string = $_ERRORS[$key];
	// }

	// return $htmlentities ? Tools::htmlentitiesUTF8(stripslashes($string)) : $string;
	return 'bbb'
}

pub fn (t Tool) get_value(error string) string {
	// global $_ERRORS;

	// if (is_null($context)) {
	// 		$context = Context::getContext();
	// }

	// @include_once(_PS_TRANSLATIONS_DIR_.$context->language->iso_code.'/errors.php');

	// if (defined('_PS_MODE_DEV_') && _PS_MODE_DEV_ && $string == 'Fatal error') {
	// 		return ('<pre>'.print_r(debug_backtrace(), true).'</pre>');
	// }

	// $key = md5(str_replace('\'', '\\\'', $string));
	// if (isset($_ERRORS)
	// 		&& is_array($_ERRORS)
	// 		&& array_key_exists($key, $_ERRORS)
	// 		&& $_ERRORS[$key] !== '') {
	// 		$string = $_ERRORS[$key];
	// }

	// return $htmlentities ? Tools::htmlentitiesUTF8(stripslashes($string)) : $string;
	return 'ssss'
}

pub fn (t Tool) get_remote_ip() string {
	// global $_ERRORS;

	// if (is_null($context)) {
	// 		$context = Context::getContext();
	// }

	// @include_once(_PS_TRANSLATIONS_DIR_.$context->language->iso_code.'/errors.php');

	// if (defined('_PS_MODE_DEV_') && _PS_MODE_DEV_ && $string == 'Fatal error') {
	// 		return ('<pre>'.print_r(debug_backtrace(), true).'</pre>');
	// }

	// $key = md5(str_replace('\'', '\\\'', $string));
	// if (isset($_ERRORS)
	// 		&& is_array($_ERRORS)
	// 		&& array_key_exists($key, $_ERRORS)
	// 		&& $_ERRORS[$key] !== '') {
	// 		$string = $_ERRORS[$key];
	// }

	// return $htmlentities ? Tools::htmlentitiesUTF8(stripslashes($string)) : $string;
	return 'aaa'
}
