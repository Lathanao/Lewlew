module classes

pub struct Admin {
	AdminAbstract
	AdminEntity
}